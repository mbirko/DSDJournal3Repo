library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.all;

entity watch is

	port
	(
		-- Input ports
		clk		: in  std_logic;
		speed		: in  std_logic;
		reset 	: in  std_logic;

		-- Output ports
		sec_1		: out std_logic_vector(6 downto 0);
		sec_10	: out std_logic_vector(6 downto 0);
		min_1		: out std_logic_vector(6 downto 0);
		min_10	: out std_logic_vector(6 downto 0);
		hrs_1		: out std_logic_vector(6 downto 0);
		hrs_10	: out std_logic_vector(6 downto 0)
		
	);
end watch;

architecture watch_impl of watch is
	-- signal from clockgen
	signal clkOutSignal	: std_logic;

	-- signals from overflow of sec, min and hrs
	signal cout_sec_1		: std_logic; 
	signal cout_sec_10	: std_logic; 
	signal cout_min_1 	: std_logic; 
	signal cout_min_10 	: std_logic; 
	signal cout_hrs_1 	: std_logic; 
	signal cout_hrs_10 	: std_logic; 
	-- signals for the value count of sec, min and hrs
	signal count_sec_1	: std_logic_vector(3 downto 0);
	signal count_sec_10	: std_logic_vector(3 downto 0);
	signal count_min_1	: std_logic_vector(3 downto 0);
	signal count_min_10	: std_logic_vector(3 downto 0);
	signal count_hrs_1	: std_logic_vector(3 downto 0);
	signal count_hrs_10	: std_logic_vector(3 downto 0);
	

	
begin
-- CLOCKGEN
	clockGen : entity clock_gen
		port map 
		(
			clk => clk,
			speed => speed,
			reset => reset,
			clk_out => clkOutSignal  
		);
		
-- MULTICOUNTER AND BIN2SEVEN FOR SEC 1
	multiCounter_sec_1 : entity multi_counter
		port map 
		(		
			count => count_sec_1,
			clk => clkOutSignal,
			cout => cout_sec_1,	
			mode => "00",
			reset => reset		
		);
		
	bin2sevenseg_sec_1 : entity bin2hex
		port map 
		(
			bin => count_sec_1,
			seg => sec_1
		);	
		
-- MULTICOUNTER AND BIN2SEVEN FOR SEC 10
	multiCounter_sec_10 : entity multi_counter
		port map 
		(		
			count => count_sec_10,
			clk => cout_sec_1,
			cout => cout_sec_10,	
			mode => "01",
			reset => reset		
		);
		
	bin2sevenseg_sec_10 : entity bin2hex
		port map 
		(
			bin => count_sec_10,
			seg => sec_10
		);	

-- MULTICOUNTER AND BIN2SEVEN FOR MIN 1
	multiCounter_min_1 : entity multi_counter
		port map 
		(		
			count => count_min_1,
			clk => cout_sec_10,
			cout => cout_min_1,	
			mode => "00",
			reset => reset		
		);
		
	bin2sevenseg_min_1 : entity bin2hex
		port map 
		(
			bin => count_min_1,
			seg => min_1
		);	
		
-- MULTICOUNTER AND BIN2SEVEN FOR MIN 10
	multiCounter_min_10 : entity multi_counter
		port map 
		(		
			count => count_min_10,
			clk => cout_min_1,
			cout => cout_min_10,	
			mode => "01",
			reset => reset		
		);
		
	bin2sevenseg_min_10 : entity bin2hex
		port map 
		(
			bin => count_min_10,
			seg => min_10
		);	
		
-- MULTICOUNTER AND BIN2SEVEN FOR HRS 1
	multiCounter_hrs_1 : entity multi_counter
		port map 
		(		
			count => count_hrs_1,
			clk => cout_min_10,
			cout => cout_hrs_1,	
			mode => "00",
			reset => reset	
		);
		
	bin2sevenseg_hrs_1 : entity bin2hex
		port map 
		(
			bin => count_hrs_1,
			seg => hrs_1
		);	
		
-- MULTICOUNTER AND BIN2SEVEN FOR HRS 10
	multiCounter_hrs_10 : entity multi_counter
		port map 
		(		
			count => count_hrs_10,
			clk => cout_hrs_1,
			cout => cout_hrs_10,	
			mode => "10",
			reset => reset		
		);
		
	bin2sevenseg_hrs_10 : entity bin2hex
		port map 
		(
			bin => count_hrs_10,
			seg => hrs_10
		);	
-- RESET LOGIC
	resetProcess : process(count_hrs_1, count_hrs_10)
	variable reset_out : integer;
	begin
		if	count_hrs_10 = "0010" then
			if count_hrs_1 = "0100" then
				reset_out := '0';
			else 
				reset_out := '1';
			end if;
		end if;
		reset => reset_out;
	end process resetProcess;
end watch_impl;

