library ieee;
use ieee.std_logic_1164.all;
use work.all;

entity nand8_tester is
	port
	(
		-- Input ports
		SW	: in  std_logic_vector(7 downto 0);

		-- Output ports
		LEDR	: out std_logic;
		
	);
end nand8_tester;

architecture nand8_impl_tester of nand8_tester is

	-- Declarations (optional)

begin

	-- Process Statement (optional)

	-- Concurrent Procedure Call (optional)

	-- Concurrent Signal Assignment (optional)

	-- Conditional Signal Assignment (optional)

	-- Selected Signal Assignment (optional)

	-- Component Instantiation Statement (optional)

	-- Generate Statement (optional)

end nand8_impl_tester;
