

library ieee;
use ieee.std_logic_1164.all;

entity guess_game is
	port
	(
		inputs : in_std_logic_vector
		-- Input ports
		<name>	: in  <type>;
		<name>	: in  <type> := <default_value>;

		-- Inout ports
		<name>	: inout <type>;

		-- Output ports
		<name>	: out <type>;
		<name>	: out <type> := <default_value>
	);
end guess_game;
